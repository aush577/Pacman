//Rom with all the walls (16x24 grid)
module mazeWalls (
						output [383:0] wallData
					  );
	
	logic [383:0] walls = 
	'{
		//maze
		1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,
		1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,
		1,0,1,1,0,1,1,0,0,1,1,0,1,1,0,1,
		1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,
		1,0,0,1,0,1,1,1,1,1,1,0,1,0,0,1,
		1,1,0,1,0,0,0,1,1,0,0,0,1,0,1,1,
		1,0,0,0,0,0,0,1,1,0,0,0,0,0,0,1,
		1,0,0,1,1,1,0,0,0,0,1,1,1,0,0,1,
		1,0,0,0,1,0,0,1,1,0,0,1,0,0,0,1,
		1,0,1,0,0,0,0,0,0,0,0,0,0,1,0,1,
		1,0,1,0,1,1,1,1,1,1,1,1,0,1,0,1,
		1,0,1,0,1,0,0,0,0,0,0,1,0,1,0,1,
		1,0,1,0,1,1,1,1,1,1,1,1,0,1,0,1,
		1,0,1,0,0,0,0,0,0,0,0,0,0,1,0,1,
		1,0,0,0,0,1,1,1,1,1,1,0,0,0,0,1,
		1,1,0,0,0,0,0,1,1,0,0,0,0,0,1,1,
		1,0,0,1,1,1,0,1,1,0,1,1,1,0,0,1,
		1,0,0,0,1,0,0,0,0,0,0,1,0,0,0,1,
		1,0,0,0,0,0,1,0,0,1,0,0,0,0,0,1,
		1,0,0,1,0,1,0,0,0,0,1,0,1,0,0,1,
		1,0,1,1,0,0,0,1,1,0,0,0,1,1,0,1,
		1,0,0,1,0,1,1,1,1,1,1,0,1,0,0,1,
		1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,
		1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1
	
	};
	
	assign wallData = walls;
	
endmodule



//module mazeWalls (
//						input [4:0] addr,
//						output [15:0] data
//					  );
//	
//	//5 addr bits = 32 spots
//	//16x24 blocks
//	logic [23:0][15:0] ROM = 
//	{
//		//maze
//		16'b 1111111111111111,
//		16'b 1000000000000001,
//		16'b 1011011001101101,
//		16'b 1000000000000001,
//		16'b 1001011111101001,
//		16'b 1101000110001011,
//		16'b 1000000110000001,
//		16'b 1001110000111001,
//		16'b 1000100110010001,
//		16'b 1010000000000101,
//		16'b 1010111111110101,
//		16'b 1010100000010101,
//		16'b 1010111001110101,
//		16'b 1010000000000101,
//		16'b 1000011111100001,
//		16'b 1100000110000011,
//		16'b 1001110110111001,
//		16'b 1000100000010001,
//		16'b 1000001001000001,
//		16'b 1001010000101001,
//		16'b 1011000110001101,
//		16'b 1001011111101001,
//		16'b 1000000000000001,
//		16'b 1111111111111111
//	
//	};
//
//	assign data = ROM[addr];
//
//
//endmodule


