module ghostSprite (
							input [6:0] addr,
							output [15:0] data
						 );
	
	//7 addr bits = 128 spots
	logic [127:0][15:0] ROM = 
	{
		//ghost
//		16'b 0000000000000000,
//		16'b 0000000000000000,
//		16'b 0000011111100000,
//		16'b 0000111111110000,
//		16'b 0001111111111000,
//		16'b 0011100110011100,
//		16'b 0011000110001100,
//		16'b 0011000110001100,
//		16'b 0011100110011100,
//		16'b 0011111111111100,
//		16'b 0011111111111100,
//		16'b 0011111111111100,
//		16'b 0011101111011100,
//		16'b 0001000110001000,
//		16'b 0000000000000000,
//		16'b 0000000000000000
	
		16'b 0000000000000000,
		16'b 0000000000000000,
		16'b 0001000110001000,
		16'b 0011101111011100,
		16'b 0011111111111100,
		16'b 0011111111111100,
		16'b 0011111111111100,
		16'b 0011100110011100,
		16'b 0011000110001100,
		16'b 0011000110001100,
		16'b 0011100110011100,
		16'b 0001111111111000,
		16'b 0000111111110000,
		16'b 0000011111100000,
		16'b 0000000000000000,
		16'b 0000000000000000
	
	};

	assign data = ROM[addr];


endmodule
