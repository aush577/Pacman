module sprites (
						input [6:0] addr,
						output [15:0] data
					);
	
	//7 addr bits = 128 spots
	logic [127:0][15:0] ROM = 
	{

		//down
		16'b 0000000000000000,
		16'b 0000000000000000,
		16'b 0000001111000000,
		16'b 0000011111100000,
		16'b 0000111111110000,
		16'b 0001111111111000,
		16'b 0011111111111100,
		16'b 0011111111111100,
		16'b 0011111111111100,
		16'b 0011111111111100,
		16'b 0001111001111000,
		16'b 0000110000110000,
		16'b 0000010000100000,
		16'b 0000000000000000,
		16'b 0000000000000000,
		16'b 0000000000000000,
		
		//up
		16'b 0000000000000000,
		16'b 0000000000000000,
		16'b 0000000000000000,
		16'b 0000010000100000,
		16'b 0000110000110000,
		16'b 0001111001111000,
		16'b 0011111111111100,
		16'b 0011111111111100,
		16'b 0011111111111100,
		16'b 0011111111111100,
		16'b 0001111111111000,
		16'b 0000111111110000,
		16'b 0000011111100000,
		16'b 0000001111000000,
		16'b 0000000000000000,
		16'b 0000000000000000,
		
		//right
		16'b 0000000000000000,
		16'b 0000000000000000,
		16'b 0000001111000000,
		16'b 0000011111100000,
		16'b 0000111111110000,
		16'b 0001111111111000,
		16'b 0011111111100000,
		16'b 0011111111000000,
		16'b 0011111111000000,
		16'b 0011111111100000,
		16'b 0001111111111000,
		16'b 0000111111110000,
		16'b 0000011111100000,
		16'b 0000001111000000,
		16'b 0000000000000000,
		16'b 0000000000000000,
		
		//left
		16'b 0000000000000000,
		16'b 0000000000000000,
		16'b 0000001111000000,
		16'b 0000011111100000,
		16'b 0000111111110000,
		16'b 0001111111111000,
		16'b 0000011111111100,
		16'b 0000001111111100,
		16'b 0000001111111100,
		16'b 0000011111111100,
		16'b 0001111111111000,
		16'b 0000111111110000,
		16'b 0000011111100000,
		16'b 0000001111000000,
		16'b 0000000000000000,
		16'b 0000000000000000
		
	
	
	};

	assign data = ROM[addr];


endmodule
