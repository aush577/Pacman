module scoreChars (
					input [3:0] addr,
					output [47:0] data
				);
	
	logic [15:0][47:0] ROM = 
	{
		// score:
		
//		48'b000000000000000000000000000000000000000000000000, 
//		48'b000000000000000000000000000000000000000000000000,
//		48'b000000000000000000000000000000000000000000000000,
//		48'b001111100001111000111110011100110111111100000000,
//		48'b011000110011001101100011001100110011001100001100,
//		48'b011000110110000101100011001100110011000100001100,
//		48'b000000110110000001100011001100110011000000000000,
//		48'b000001100110000001100011001101100011010000000000,
//		48'b000111000110000001100011001111100011110000000000,
//		48'b001100000110000001100011001100110011010000001100,
//		48'b011000110110000101100011001100110011000100001100,
//		48'b011000110011001101100011001100110011001100000000,
//		48'b001111100001111000111110011111100111111100000000,
//		48'b000000000000000000000000000000000000000000000000,
//		48'b000000000000000000000000000000000000000000000000,
//		48'b000000000000000000000000000000000000000000000000   
		
		
		48'b000000000000000000000000000000000000000000000000,
		48'b000000000000000000000000000000000000000000000000,
		48'b000000000000000000000000000000000000000000000000,
		48'b000000000000000000000000000000000000000000000000,
		48'b000000000000000000000000000000000000000000000000,
		48'b000000001111111011001110011111000111100001111100,
		48'b001100001100110011001100110001101100110011000110,
		48'b001100001000110011001100110001101000011011000110,
		48'b000000000000110011001100110001100000011011000000,
		48'b000000000010110001101100110001100000011001100000,
		48'b000000000011110001111100110001100000011000111000,
		48'b001100000010110011001100110001100000011000001100,
		48'b001100001000110011001100110001101000011011000110,
		48'b000000001100110011001100110001101100110011000110,
		48'b000000001111111001111110011111000111100001111100,
		48'b000000000000000000000000000000000000000000000000

		
		
//		48'b000000000000000000000000000000000000000000000000,   
//		48'b000000000000000000000000000000000000000000000000,
//		48'b000000000000000000000000000000000000000000000000,
//		48'b001111100001111000111110011111100111111100000000,
//		48'b011000110011001101100011001100110011001100000000,
//		48'b011000110110000101100011001100110011000100001100,
//		48'b001100000110000001100011001100110011010000001100,
//		48'b000111000110000001100011001111100011110000000000,
//		48'b000001100110000001100011001101100011010000000000,
//		48'b000000110110000001100011001100110011000000000000,
//		48'b011000110110000101100011001100110011000100001100,
//		48'b011000110011001101100011001100110011001100001100,
//		48'b001111100001111000111110011100110111111100000000,
//		48'b000000000000000000000000000000000000000000000000,
//		48'b000000000000000000000000000000000000000000000000,
//		48'b000000000000000000000000000000000000000000000000                    
	};
	
	assign data = ROM[addr];

endmodule 