module maze (
					input [8:0] addr,
					output [255:0] data
				);
	
	//9 addr bits = 512 spots
	//16x24 (16 bit blocks) maze = 256x384
	//16 bit blocks = 0000 or ffff
	//Reverse addresses for y axis counter
	logic [511:0][255:0] ROM = 
	{
	
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111,
			256'b 1111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111,
			256'b 1111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111,
			256'b 1111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111,
			256'b 1111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111,
			256'b 1111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111,
			256'b 1111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111,
			256'b 1111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111,
			256'b 1111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111,
			256'b 1111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111,
			256'b 1111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111,
			256'b 1111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111,
			256'b 1111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111,
			256'b 1111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111,
			256'b 1111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111,
			256'b 1111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111,
			256'b 1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111,
			256'b 1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111,
			256'b 1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111,
			256'b 1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111,
			256'b 1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111,
			256'b 1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111,
			256'b 1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111,
			256'b 1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111,
			256'b 1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111,
			256'b 1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111,
			256'b 1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111,
			256'b 1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111,
			256'b 1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111,
			256'b 1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111,
			256'b 1111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000111111111111111111111111111111110000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000001111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111,
			256'b 1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111

	
	};


	assign data = ROM[addr];


endmodule
