module numbers (
					input [7:0] addr,
					output [7:0] data
				);
	
	logic [255:0][7:0] ROM = 
	{
	
		8'b00000000,
		8'b00000000,
		8'b00000000,
		8'b00000000,
		8'b00011110,
		8'b00110000,
		8'b01100000,
		8'b01100000,
		8'b01100000,
		8'b01111110,
		8'b01100011,
		8'b01100011,
		8'b01100011,
		8'b00111110,
		8'b00000000,
		8'b00000000,

		8'b00000000,
		8'b00000000,
		8'b00000000,
		8'b00000000,
		8'b00111110,
		8'b01100011,
		8'b01100011,
		8'b01100011,
		8'b01100011,
		8'b00111110,
		8'b01100011,
		8'b01100011,
		8'b01100011,
		8'b00111110,
		8'b00000000,
		8'b00000000,

		8'b00000000,
		8'b00000000,
		8'b00000000,
		8'b00000000,
		8'b00001100,
		8'b00001100,
		8'b00001100,
		8'b00001100,
		8'b00011000,
		8'b00110000,
		8'b01100000,
		8'b01100000,
		8'b01100011,
		8'b01111111,
		8'b00000000,
		8'b00000000,

		8'b00000000,
		8'b00000000,
		8'b00000000,
		8'b00000000,
		8'b00111110,
		8'b01100011,
		8'b01100011,
		8'b01100011,
		8'b01100011,
		8'b00111111,
		8'b00000011,
		8'b00000011,
		8'b00000110,
		8'b00011100,
		8'b00000000,
		8'b00000000,

		8'b00000000,
		8'b00000000,
		8'b00000000,
		8'b00000000,
		8'b00111110,
		8'b01100011,
		8'b01100000,
		8'b01100000,
		8'b01100000,
		8'b00111111,
		8'b00000011,
		8'b00000011,
		8'b00000011,
		8'b01111111,
		8'b00000000,
		8'b00000000,

		8'b00000000,
		8'b00000000,
		8'b00000000,
		8'b00000000,
		8'b01111000,
		8'b00110000,
		8'b00110000,
		8'b00110000,
		8'b01111111,
		8'b00110011,
		8'b00110110,
		8'b00111100,
		8'b00111000,
		8'b00110000,
		8'b00000000,
		8'b00000000,

		8'b00000000,
		8'b00000000,
		8'b00000000,
		8'b00000000,
		8'b00111110,
		8'b01100011,
		8'b01100000,
		8'b01100000,
		8'b01100000,
		8'b00111100,
		8'b01100000,
		8'b01100000,
		8'b01100011,
		8'b00111110,
		8'b00000000,
		8'b00000000,

		8'b00000000,
		8'b00000000,
		8'b00000000,
		8'b00000000,
		8'b01111111,
		8'b01100011,
		8'b00000011,
		8'b00000110,
		8'b00001100,
		8'b00011000,
		8'b00110000,
		8'b01100000,
		8'b01100011,
		8'b00111110,
		8'b00000000,
		8'b00000000,

		8'b00000000,
		8'b00000000,
		8'b00000000,
		8'b00000000,
		8'b01111110,
		8'b00011000,
		8'b00011000,
		8'b00011000,
		8'b00011000,
		8'b00011000,
		8'b00011000,
		8'b00011110,
		8'b00011100,
		8'b00011000,
		8'b00000000,
		8'b00000000,

		8'b00000000,
		8'b00000000,
		8'b00000000,
		8'b00000000,
		8'b00111110,
		8'b01100011,
		8'b01100011,
		8'b01100111,
		8'b01101111,
		8'b01111011,
		8'b01110011,
		8'b01100011,
		8'b01100011,
		8'b00111110,
		8'b00000000

		
		
	
	
	
//		8'b00000000, // 0
//		8'b00000000, // 1
//		8'b01111100, // 2  *****
//		8'b11000110, // 3 **   **
//		8'b11000110, // 4 **   **
//		8'b11000110, // 5 **   **
//		8'b01111110, // 6  ******
//		8'b00000110, // 7      **
//		8'b00000110, // 8      **
//		8'b00000110, // 9      **
//		8'b00001100, // a     **
//		8'b01111000, // b  ****
//		8'b00000000, // c
//		8'b00000000, // d
//		8'b00000000, // e
//		8'b00000000, // f
//
//		8'b00000000, // 0
//		8'b00000000, // 1
//		8'b01111100, // 2  *****
//		8'b11000110, // 3 **   **
//		8'b11000110, // 4 **   **
//		8'b11000110, // 5 **   **
//		8'b01111100, // 6  *****
//		8'b11000110, // 7 **   **
//		8'b11000110, // 8 **   **
//		8'b11000110, // 9 **   **
//		8'b11000110, // a **   **
//		8'b01111100, // b  *****
//		8'b00000000, // c
//		8'b00000000, // d
//		8'b00000000, // e
//		8'b00000000, // f
//	
//		8'b00000000, // 0
//		8'b00000000, // 1
//		8'b11111110, // 2 *******
//		8'b11000110, // 3 **   **
//		8'b00000110, // 4      **
//		8'b00000110, // 5      **
//		8'b00001100, // 6     **
//		8'b00011000, // 7    **
//		8'b00110000, // 8   **
//		8'b00110000, // 9   **
//		8'b00110000, // a   **
//		8'b00110000, // b   **
//		8'b00000000, // c
//		8'b00000000, // d
//		8'b00000000, // e
//		8'b00000000, // f
//
//		8'b00000000, // 0
//		8'b00000000, // 1
//		8'b00111000, // 2   ***
//		8'b01100000, // 3  **
//		8'b11000000, // 4 **
//		8'b11000000, // 5 **
//		8'b11111100, // 6 ******
//		8'b11000110, // 7 **   **
//		8'b11000110, // 8 **   **
//		8'b11000110, // 9 **   **
//		8'b11000110, // a **   **
//		8'b01111100, // b  *****
//		8'b00000000, // c
//		8'b00000000, // d
//		8'b00000000, // e
//		8'b00000000, // f
//
//		8'b00000000, // 0
//		8'b00000000, // 1
//		8'b11111110, // 2 *******
//		8'b11000000, // 3 **
//		8'b11000000, // 4 **
//		8'b11000000, // 5 **
//		8'b11111100, // 6 ******
//		8'b00000110, // 7      **
//		8'b00000110, // 8      **
//		8'b00000110, // 9      **
//		8'b11000110, // a **   **
//		8'b01111100, // b  *****
//		8'b00000000, // c
//		8'b00000000, // d
//		8'b00000000, // e
//		8'b00000000, // f
//
//		8'b00000000, // 0
//		8'b00000000, // 1
//		8'b00001100, // 2     **
//		8'b00011100, // 3    ***
//		8'b00111100, // 4   ****
//		8'b01101100, // 5  ** **
//		8'b11001100, // 6 **  **
//		8'b11111110, // 7 *******
//		8'b00001100, // 8     **
//		8'b00001100, // 9     **
//		8'b00001100, // a     **
//		8'b00011110, // b    ****
//		8'b00000000, // c
//		8'b00000000, // d
//		8'b00000000, // e
//		8'b00000000, // f
//
//		8'b00000000, // 0
//		8'b00000000, // 1
//		8'b01111100, // 2  *****
//		8'b11000110, // 3 **   **
//		8'b00000110, // 4      **
//		8'b00000110, // 5      **
//		8'b00111100, // 6   ****
//		8'b00000110, // 7      **
//		8'b00000110, // 8      **
//		8'b00000110, // 9      **
//		8'b11000110, // a **   **
//		8'b01111100, // b  *****
//		8'b00000000, // c
//		8'b00000000, // d
//		8'b00000000, // e
//		8'b00000000, // f
//
//		8'b00000000, // 0
//		8'b00000000, // 1
//		8'b01111100, // 2  *****
//		8'b11000110, // 3 **   **
//		8'b00000110, // 4      **
//		8'b00001100, // 5     **
//		8'b00011000, // 6    **
//		8'b00110000, // 7   **
//		8'b01100000, // 8  **
//		8'b11000000, // 9 **
//		8'b11000110, // a **   **
//		8'b11111110, // b *******
//		8'b00000000, // c
//		8'b00000000, // d
//		8'b00000000, // e
//		8'b00000000, // f
//
//		8'b00000000, // 0
//		8'b00000000, // 1
//		8'b00011000, // 2
//		8'b00111000, // 3
//		8'b01111000, // 4    **
//		8'b00011000, // 5   ***
//		8'b00011000, // 6  ****
//		8'b00011000, // 7    **
//		8'b00011000, // 8    **
//		8'b00011000, // 9    **
//		8'b00011000, // a    **
//		8'b01111110, // b    **
//		8'b00000000, // c    **
//		8'b00000000, // d  ******
//		8'b00000000, // e
//		8'b00000000, // f
//
//		8'b00000000, // 0
//		8'b00000000, // 1
//		8'b01111100, // 2  *****
//		8'b11000110, // 3 **   **
//		8'b11000110, // 4 **   **
//		8'b11001110, // 5 **  ***
//		8'b11011110, // 6 ** ****
//		8'b11110110, // 7 **** **
//		8'b11100110, // 8 ***  **
//		8'b11000110, // 9 **   **
//		8'b11000110, // a **   **
//		8'b01111100, // b  *****
//		8'b00000000, // c
//		8'b00000000, // d
//		8'b00000000, // e
//		8'b00000000 // f



	
	
	
//			// code x0
//		8'b00000000, // 0
//		8'b00000000, // 1
//		8'b01111100, // 2  *****
//		8'b11000110, // 3 **   **
//		8'b11000110, // 4 **   **
//		8'b11001110, // 5 **  ***
//		8'b11011110, // 6 ** ****
//		8'b11110110, // 7 **** **
//		8'b11100110, // 8 ***  **
//		8'b11000110, // 9 **   **
//		8'b11000110, // a **   **
//		8'b01111100, // b  *****
//		8'b00000000, // c
//		8'b00000000, // d
//		8'b00000000, // e
//		8'b00000000, // f
//		// code x16
//		8'b00000000, // 0
//		8'b00000000, // 1
//		8'b00011000, // 2
//		8'b00111000, // 3
//		8'b01111000, // 4    **
//		8'b00011000, // 5   ***
//		8'b00011000, // 6  ****
//		8'b00011000, // 7    **
//		8'b00011000, // 8    **
//		8'b00011000, // 9    **
//		8'b00011000, // a    **
//		8'b01111110, // b    **
//		8'b00000000, // c    **
//		8'b00000000, // d  ******
//		8'b00000000, // e
//		8'b00000000, // f
//		// code x32
//		8'b00000000, // 0
//		8'b00000000, // 1
//		8'b01111100, // 2  *****
//		8'b11000110, // 3 **   **
//		8'b00000110, // 4      **
//		8'b00001100, // 5     **
//		8'b00011000, // 6    **
//		8'b00110000, // 7   **
//		8'b01100000, // 8  **
//		8'b11000000, // 9 **
//		8'b11000110, // a **   **
//		8'b11111110, // b *******
//		8'b00000000, // c
//		8'b00000000, // d
//		8'b00000000, // e
//		8'b00000000, // f
//		// code x33
//		8'b00000000, // 0
//		8'b00000000, // 1
//		8'b01111100, // 2  *****
//		8'b11000110, // 3 **   **
//		8'b00000110, // 4      **
//		8'b00000110, // 5      **
//		8'b00111100, // 6   ****
//		8'b00000110, // 7      **
//		8'b00000110, // 8      **
//		8'b00000110, // 9      **
//		8'b11000110, // a **   **
//		8'b01111100, // b  *****
//		8'b00000000, // c
//		8'b00000000, // d
//		8'b00000000, // e
//		8'b00000000, // f
//		// code x34
//		8'b00000000, // 0
//		8'b00000000, // 1
//		8'b00001100, // 2     **
//		8'b00011100, // 3    ***
//		8'b00111100, // 4   ****
//		8'b01101100, // 5  ** **
//		8'b11001100, // 6 **  **
//		8'b11111110, // 7 *******
//		8'b00001100, // 8     **
//		8'b00001100, // 9     **
//		8'b00001100, // a     **
//		8'b00011110, // b    ****
//		8'b00000000, // c
//		8'b00000000, // d
//		8'b00000000, // e
//		8'b00000000, // f
//		// code x35
//		8'b00000000, // 0
//		8'b00000000, // 1
//		8'b11111110, // 2 *******
//		8'b11000000, // 3 **
//		8'b11000000, // 4 **
//		8'b11000000, // 5 **
//		8'b11111100, // 6 ******
//		8'b00000110, // 7      **
//		8'b00000110, // 8      **
//		8'b00000110, // 9      **
//		8'b11000110, // a **   **
//		8'b01111100, // b  *****
//		8'b00000000, // c
//		8'b00000000, // d
//		8'b00000000, // e
//		8'b00000000, // f
//		// code x36
//		8'b00000000, // 0
//		8'b00000000, // 1
//		8'b00111000, // 2   ***
//		8'b01100000, // 3  **
//		8'b11000000, // 4 **
//		8'b11000000, // 5 **
//		8'b11111100, // 6 ******
//		8'b11000110, // 7 **   **
//		8'b11000110, // 8 **   **
//		8'b11000110, // 9 **   **
//		8'b11000110, // a **   **
//		8'b01111100, // b  *****
//		8'b00000000, // c
//		8'b00000000, // d
//		8'b00000000, // e
//		8'b00000000, // f
//		// code x37
//		8'b00000000, // 0
//		8'b00000000, // 1
//		8'b11111110, // 2 *******
//		8'b11000110, // 3 **   **
//		8'b00000110, // 4      **
//		8'b00000110, // 5      **
//		8'b00001100, // 6     **
//		8'b00011000, // 7    **
//		8'b00110000, // 8   **
//		8'b00110000, // 9   **
//		8'b00110000, // a   **
//		8'b00110000, // b   **
//		8'b00000000, // c
//		8'b00000000, // d
//		8'b00000000, // e
//		8'b00000000, // f
//		// code x38
//		8'b00000000, // 0
//		8'b00000000, // 1
//		8'b01111100, // 2  *****
//		8'b11000110, // 3 **   **
//		8'b11000110, // 4 **   **
//		8'b11000110, // 5 **   **
//		8'b01111100, // 6  *****
//		8'b11000110, // 7 **   **
//		8'b11000110, // 8 **   **
//		8'b11000110, // 9 **   **
//		8'b11000110, // a **   **
//		8'b01111100, // b  *****
//		8'b00000000, // c
//		8'b00000000, // d
//		8'b00000000, // e
//		8'b00000000, // f
//		// code x39
//		8'b00000000, // 0
//		8'b00000000, // 1
//		8'b01111100, // 2  *****
//		8'b11000110, // 3 **   **
//		8'b11000110, // 4 **   **
//		8'b11000110, // 5 **   **
//		8'b01111110, // 6  ******
//		8'b00000110, // 7      **
//		8'b00000110, // 8      **
//		8'b00000110, // 9      **
//		8'b00001100, // a     **
//		8'b01111000, // b  ****
//		8'b00000000, // c
//		8'b00000000, // d
//		8'b00000000, // e
//		8'b00000000 // f
	};
	
	assign data = ROM[addr];

endmodule 