module gameOver(
					input [3:0] addr,
					output [71:0] data
				);

	logic [15:0][71:0] ROM =
	{
	
		72'b000000000000000000000000000000000000000000000000000000000000000000000000,
		72'b000000000000000000000000000000000000000000000000000000000000000000000000,
		72'b000000000000000000000000000000000000000000000000000000000000000000000000,
		72'b011001110111111100011000001111100000000001111111110000110110001101011100,
		72'b011001100110011000111100011000110000000001100110110000110110001101100110,
		72'b011001100100011001100110011000110000000001000110110000110110001101100011,
		72'b011001100000011011000011011000110000000000000110110000110110001101100011,
		72'b001101100001011011000011011000110000000000010110110000110111111101111011,
		72'b001111100001111011000011011000110000000000011110110110110110001100000011,
		72'b011001100001011011000011011000110000000000010110111111110110001100000011,
		72'b011001100100011011000011011000110000000001000110111111110011011001000011,
		72'b011001100110011011000011011000110000000001100110111001110001110001100110,
		72'b001111110111111111000011001111100000000001111111110000110000100000111100,
		72'b000000000000000000000000000000000000000000000000000000000000000000000000,
		72'b000000000000000000000000000000000000000000000000000000000000000000000000,
		72'b000000000000000000000000000000000000000000000000000000000000000000000000




	
	
//		72'b000000000000000000000000000000000000000000000000000000000000000000000000,
//		72'b000000000000000000000000000000000000000000000000000000000000000000000000,
//		72'b000000000000000000000000000000000000000000000000000000000000000000000000,
//		72'b001111000001000011000011111111100000000001111100110000111111111011111100,
//		72'b011001100011100011100111011001100000000011000110110000110110011001100110,
//		72'b110000100110110011111111011000100000000011000110110000110110001001100110,
//		72'b110000001100011011111111011010000000000011000110110000110110100001100110,
//		72'b110000001100011011011011011110000000000011000110110000110111100001111100,
//		72'b110111101111111011000011011010000000000011000110110000110110100001101100,
//		72'b110001101100011011000011011000000000000011000110110000110110000001100110,
//		72'b110001101100011011000011011000100000000011000110011001100110001001100110,
//		72'b011001101100011011000011011001100000000011000110001111000110011001100110,
//		72'b001110101100011011000011111111100000000001111100000110001111111011100110,
//		72'b000000000000000000000000000000000000000000000000000000000000000000000000,
//		72'b000000000000000000000000000000000000000000000000000000000000000000000000,
//		72'b000000000000000000000000000000000000000000000000000000000000000000000000
	};

assign data = ROM[addr];

endmodule
